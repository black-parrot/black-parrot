
package bp_fe_icache_pkg;

`include "bp_common_lce_cce_if.vh"
`include "bsg_defines.v"

endpackage : bp_fe_icache_pkg
