/*
 * bp_me_pkg.vh
 *
 * Contains the interface structures used for communicating between the CCE and Memory.
 *
 */

package bp_me_pkg;

  `include "bsg_defines.v"
  `include "bp_common_mem_if.vh"

endpackage : bp_me_pkg

