package itlb_pkg;

localparam bp_ppn_width_gp = 44;
localparam bp_ppn_start_bit_gp = 12;
endpackage : itlb_pkg
