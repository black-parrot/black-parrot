
module bp_be_nonsynth_dcache_tracer
 import bp_common_pkg::*;
 import bp_common_aviary_pkg::*;
 import bp_be_pkg::*;
 import bp_common_rv64_pkg::*;
 #(parameter bp_params_e bp_params_p = e_bp_inv_cfg
   `declare_bp_proc_params(bp_params_p)
   `declare_bp_cache_service_if_widths(paddr_width_p, ptag_width_p, lce_sets_p, dcache_assoc_p, dword_width_p, cce_block_width_p, dcache)
   
   // Default parameters
   , parameter dcache_trace_file_p = "dcache"

   // Calculated parameters
   , localparam mhartid_width_lp      = `BSG_SAFE_CLOG2(num_core_p)
   , localparam block_size_in_words_lp=dcache_assoc_p
   , localparam cache_block_multiplier_width_lp = 2**(3-`BSG_SAFE_CLOG2(dcache_assoc_p))
   , localparam cache_block_width_lp = dword_width_p * cache_block_multiplier_width_lp
   , localparam data_mem_mask_width_lp=(cache_block_width_lp>>3)
   , localparam bypass_data_width_lp = (dword_width_p >> 3)
   , localparam byte_offset_width_lp=`BSG_SAFE_CLOG2(cache_block_width_lp>>3)
   , localparam word_offset_width_lp=`BSG_SAFE_CLOG2(block_size_in_words_lp)
   , localparam block_offset_width_lp=(word_offset_width_lp+byte_offset_width_lp)
   , localparam index_width_lp=`BSG_SAFE_CLOG2(lce_sets_p)
   , localparam ptag_width_lp=(paddr_width_p-bp_page_offset_width_gp)
   , localparam way_id_width_lp=`BSG_SAFE_CLOG2(dcache_assoc_p)
  
   , localparam lce_data_width_lp=(lce_assoc_p*dword_width_p)

   )
  (  input                                                 clk_i
   , input                                                 reset_i
   , input                                                 freeze_i
   , input [mhartid_width_lp-1:0]                          mhartid_i
      
   // Tag lookup
   , input                                                 v_tl_r
   
   // Tag Verify
   , input                                                 v_tv_r
   , input [paddr_width_p-1:0]                             paddr_tv_r
   , input                                                 lr_miss_tv
   , input                                                 sc_op_tv_r
   , input                                                 sc_success

   // Miss Packet
   , input                                                 cache_req_v_o
   , input [dcache_req_width_lp-1:0]                       cache_req_o

   // Cache Metadata
   , input [dcache_req_metadata_width_lp-1:0]              cache_req_metadata_o 
   , input                                                 cache_req_metadata_v_o

   , input                                                 cache_req_complete_i

   // Cache data
   , input                                                 v_o
   , input [dword_width_p-1:0]                             load_data
   , input                                                 dcache_miss_o
   , input [dword_width_p-1:0]                             store_data

   // Fill Packets
   , input                                                 data_mem_pkt_v_i
   , input [dcache_data_mem_pkt_width_lp-1:0]              data_mem_pkt_i
   , input                                                 data_mem_pkt_ready_o

   , input                                                 tag_mem_pkt_v_i
   , input [dcache_tag_mem_pkt_width_lp-1:0]               tag_mem_pkt_i
   , input                                                 tag_mem_pkt_ready_o

   , input                                                 stat_mem_pkt_v_i
   , input [dcache_stat_mem_pkt_width_lp-1:0]              stat_mem_pkt_i
   , input                                                 stat_mem_pkt_ready_o
   );

  `declare_bp_cache_service_if(paddr_width_p, ptag_width_p, lce_sets_p, dcache_assoc_p, dword_width_p, cce_block_width_p, dcache);

  // Input Casting  
  bp_dcache_req_s cache_req_cast_o;
  bp_dcache_req_metadata_s cache_req_metadata_cast_o;
  assign cache_req_cast_o = cache_req_o;
  assign cache_req_metadata_cast_o = cache_req_metadata_o;

  bp_dcache_data_mem_pkt_s data_mem_pkt_cast_i;
  bp_dcache_tag_mem_pkt_s tag_mem_pkt_cast_i;
  bp_dcache_stat_mem_pkt_s stat_mem_pkt_cast_i;
  assign data_mem_pkt_cast_i = data_mem_pkt_i; 
  assign tag_mem_pkt_cast_i = tag_mem_pkt_i;
  assign stat_mem_pkt_cast_i = stat_mem_pkt_i;

  integer file;
  string file_name;
  
  wire delay_li = reset_i | freeze_i;
  always_ff @(negedge delay_li)
   begin
     file_name = $sformatf("%s_%x.trace", dcache_trace_file_p, mhartid_i);
     file      = $fopen(file_name, "w");
   end

  string op;

  always_comb begin
      if (lr_miss_tv & cache_req_v_o)
        op = "[lr]";
      else if(sc_op_tv_r)
        op = "[sc]";
      else if (cache_req_v_o & cache_req_cast_o.msg_type == e_miss_store)
        op = "[store]";
      else if (cache_req_v_o & cache_req_cast_o.msg_type == e_miss_load)
        op = "[load]";
      else if (cache_req_v_o & cache_req_cast_o.msg_type == e_uc_load)
        op = "[uncached load]";
      else if (cache_req_v_o & cache_req_cast_o.msg_type == e_uc_store)
        op = "[uncached store]";
      else if (cache_req_v_o & cache_req_cast_o.msg_type == e_cache_flush)
        op = "[fencei req]";
      else
        op = "[null]";
    end

  always_ff @(posedge clk_i) begin
 
      if(v_tl_r) 
        $fwrite(file, "[%t] tag_lookup: %x \n", $time, v_tl_r);
      
      if(v_tv_r)
        $fwrite(file, "[%t] tag_verify: %x \n", $time, v_tv_r);
      
      if(sc_success)
        $fwrite(file, "SC SUCEESS! \n");
      
      
      if (cache_req_v_o) begin
        $fwrite(file, "[%t] valid cache_req: %x \n", $time, cache_req_v_o);
        $fwrite(file, "[%t] %s addr: %x data: %x cache_miss: %x \n", $time, op, cache_req_cast_o.addr, cache_req_cast_o.data, dcache_miss_o);
      end

      if (cache_req_metadata_v_o)
        $fwrite(file, "[%t] lru_way: %x dirty: %x \n", $time, cache_req_metadata_cast_o.repl_way, cache_req_metadata_cast_o.dirty);
      
      if (cache_req_complete_i)
        $fwrite(file, "[%t] Cache request completed \n", $time);

      if (data_mem_pkt_v_i)
        $fwrite(file, "[%t] Data Mem: op: %x index: %x data: %x \n", $time, data_mem_pkt_cast_i.opcode, data_mem_pkt_cast_i.index, data_mem_pkt_cast_i.data);

      if (tag_mem_pkt_v_i)
        $fwrite(file, "[%t] Tag Mem: op: %x index: %x tag: %x state: %x \n", $time, tag_mem_pkt_cast_i.opcode, tag_mem_pkt_cast_i.index, tag_mem_pkt_cast_i.tag, tag_mem_pkt_cast_i.state);

      if (stat_mem_pkt_v_i)
        $fwrite(file, "[%t] Stat Mem: op: %x, index: %x \n", $time, stat_mem_pkt_cast_i.opcode, stat_mem_pkt_cast_i.index);

      if (v_o)
        $fwrite(file, "[%t] load data: %x \n", $time, load_data);

      if (cache_req_v_o & (cache_req_cast_o.msg_type == e_miss_store || cache_req_cast_o.msg_type == e_uc_store))
        $fwrite(file, "[%t] store data: %x \n", $time, store_data);
    end

endmodule
