/**
 *
 * Name:
 *   bp_me_nonsynth_dev_tracer.sv
 *
 * Description:
 *
 */

`include "bp_common_defines.svh"
`include "bp_me_defines.svh"

module bp_me_nonsynth_dev_tracer
  import bp_common_pkg::*;
  import bp_me_pkg::*;
  #(parameter bp_params_e bp_params_p = e_bp_default_cfg
    `declare_bp_proc_params(bp_params_p)

    , parameter trace_file_p = "dev"

    `declare_bp_bedrock_if_widths(paddr_width_p, lce_id_width_p, cce_id_width_p, did_width_p, lce_assoc_p)
  )
  (input                                            clk_i
   , input                                          reset_i

   , input [core_id_width_p-1:0]                    mhartid_i

   // CCE-MEM Interface
   // BedRock Stream protocol: ready&valid
   , input [mem_fwd_header_width_lp-1:0]            mem_fwd_header_i
   , input [bedrock_fill_width_p-1:0]               mem_fwd_data_i
   , input                                          mem_fwd_v_i
   , input                                          mem_fwd_ready_and_i

   , input [mem_rev_header_width_lp-1:0]            mem_rev_header_i
   , input [bedrock_fill_width_p-1:0]               mem_rev_data_i
   , input                                          mem_rev_v_i
   , input                                          mem_rev_ready_and_i
  );

  `declare_bp_bedrock_if(paddr_width_p, lce_id_width_p, cce_id_width_p, did_width_p, lce_assoc_p);

  `bp_cast_i(bp_bedrock_mem_fwd_header_s, mem_fwd_header);
  `bp_cast_i(bp_bedrock_mem_rev_header_s, mem_rev_header);

  integer file;
  string file_name;

  always_ff @(negedge reset_i)
    begin
      file_name = $sformatf("%s_%x.trace", trace_file_p, mhartid_i);
      file      = $fopen(file_name, "w");
    end

  // Tracer
  always_ff @(negedge clk_i) begin
    if (~reset_i) begin
      if (mem_fwd_v_i & mem_fwd_ready_and_i) begin
        $fdisplay(file, "%12t |: MEM FWD addr[%H] msg[%b] size[%b]"
                 , $time
                 , mem_fwd_header_cast_i.addr
                 , mem_fwd_header_cast_i.msg_type.fwd
                 , mem_fwd_header_cast_i.size
                 );
        if (mem_fwd_header_cast_i.msg_type.fwd == e_bedrock_mem_wr) begin
          $fdisplay(file, "%12t |: MEM FWD DATA %H"
                   , $time
                   , mem_fwd_data_i
                   );
        end
      end
      if (mem_rev_v_i & mem_rev_ready_and_i) begin
        $fdisplay(file, "%12t |: MEM REV addr[%H] msg[%b] size[%b]"
                 , $time
                 , mem_rev_header_cast_i.addr
                 , mem_rev_header_cast_i.msg_type.rev
                 , mem_rev_header_cast_i.size
                 );
        if (mem_rev_header_cast_i.msg_type.rev == e_bedrock_mem_rd) begin
          $fdisplay(file, "%12t |: MEM REV DATA %H"
                   , $time
                   , mem_rev_data_i
                   );
        end
      end
    end // reset & trace
  end // always_ff

endmodule
