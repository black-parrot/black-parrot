package pc_gen_pkg;

//localparam vaddr_width_p = 64;
//localparam paddr_width_p = 56;
//localparam asid_width_p  = 10;
//localparam branch_metadata_fwd_width_p = 64 + 9 + 5;

localparam __ERROR__MSG__ = "\033[31m\033[1m [ERROR] \033[0m ";
localparam __INFO__MSG__  = "\033[37m\033[1m [INFO] \033[0m ";
localparam __DEBUG__MSG__ = "\033[36m\033[1m [DEBUG] \033[0m ";

endpackage : pc_gen_pkg
