
  `include "bp_top_defines.svh"

package bp_top_pkg;

endpackage

