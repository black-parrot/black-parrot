/*
 * bp_me_pkg.vh
 *
 * Contains the interface structures used for communicating between the CCE and Memory.
 *
 */

package bp_me_pkg;

  `include "bsg_defines.v"
  `include "bp_me_cce_mem_if.vh"
  `include "bp_me_cce_io_if.vh"

endpackage : bp_me_pkg

