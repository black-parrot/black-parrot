/*
 * bp_me_pkg.vh
 *
 * Contains the interface structures used for communicating between the CCE and Memory.
 *
 */

package bp_me_pkg;

  `include "bsg_defines.v"
  `include "bp_common_mem_if.vh"
  `include "bp_mem_wormhole.vh"

endpackage : bp_me_pkg

