
package bp_fe_icache_pkg;

  `include "bp_common_bedrock_if.svh"
  `include "bsg_defines.v"
  `include "bp_fe_icache.svh"

endpackage

