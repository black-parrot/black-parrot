
package bp_fe_pkg;

  `include "bsg_defines.v"
  `include "bp_common_core_if.svh"
  `include "bp_fe_defines.svh"
  `include "bp_fe_mem_defines.svh"

endpackage : bp_fe_pkg
