
package bp_fe_pkg;

  `include "bsg_defines.v"
  `include "bp_common_fe_be_if.vh"
  `include "bp_fe_top.vh"
  `include "bp_fe_icache.vh"
  `include "bp_fe_mem_defines.vh"

endpackage : bp_fe_pkg
