`ifndef BP_COMMON_DEFINES_VH
`define BP_COMMON_DEFINES_VH

  `include "bsg_defines.v"
  `include "bp_common_defines.svh"
  `include "bp_common_core_if.svh"
  `include "bp_common_bedrock_if.svh"
  `include "bp_common_cache_engine_if.svh"
  `include "bp_common_cfg_bus_defines.svh"
  `include "bp_common_log_defines.svh"
  `include "bp_common_rv64_instr_defines.svh"
  `include "bp_common_rv64_csr_defines.svh"

`endif

