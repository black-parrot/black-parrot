/**
 *
 * Name:
 *   bp_me_wrap_counter.sv
 *
 * Description:
 *   This module generates a wrap-around count given an initial count and transaction size, for
 *   a fixed maximum count. Both the initial count and transaction size are zero-based.
 *   This count can be used to generate the word bits of a protocol message address.
 *
 *   max_val_p is equal to the maximum count - 1 (i.e., it is zero-based).
 *   max_val_p+1 must be a power of two for the wrap-around counting to work properly.
 *   For a protocol message, max_val_p is equal to (block width / stream width) - 1.
 *   E.g., if a block is divided into 8 words, max_val_p = 7.
 *
 *   size_i is the zero-based transaction size (e.g., a transaction of 4 words has size_i = 3).
 *   size_i+1 must be a power of two for the wrap-around count to work. If size_i+1 is not a
 *   power of two, the count wraps as if size_i+1 is the next power of two.
 *   (e.g., max_val_p = 3, then size_i = 2 wraps same as size_i = 3)
 *
 *   val_i is the zero-based initial word in [0, max_val_p] of the transaction.
 *   Both size_i and val_i must be held constant throughout the transaction.
 *
 *   en_i increments the count output on wrap_o
 *
 *   wrap_o is a count that wraps around at the end of the naturally aligned sub-block with
 *   size (size_i+1). The count is wrapped within the size_i aligned portion of [0, max_val_p]
 *   that includes val_i.
 *
 *   first_o is raised when wrap_o is the first count of the sequence.
 *   last_o is raised when wrap_o is the last count of the sequence, and depends on size_i.
 *
 *   The following describes how this wrap-around counting can be used to generate the word bits
 *   of an address. This is useful for transmitting a block of data as sequence or stream of
 *   words where (block width / stream data channel width) = max_val_p + 1.
 *
 *   A canonical block address can be viewed as:
 *   __________________________________________________________
 *   |                |          block offset                  |  block address
 *   |  upper address |________________________________________|
 *   |                |   stream count /   |  stream offset /  |  stream word address
 *   |                |   word address     |  word byte offset |
 *   |________________|____________________|___________________|
 *
 *   where stream offset is a byte offset of the current stream word and stream count is
 *   the index of the word in the block in the range [0, max_val_p]. This module computes
 *   the stream count or word address as the wrap_o output.
 *
 *   To produce wrap_o, the stream count / word address is further divided into:
 *   __________________________________________________
 *   |    sub-block number     |    sub-block count    |
 *   |_________________________|_______________________|
 *
 *   For a given sequence of wrap_o, the sub-block number portion of wrap_o remains constant
 *   while the sub-block count portion is generated by a counter. The number of bits
 *   derived from the counter versus the initial stream word input (val_i) is determined by
 *   the transaction size (size_i) input. A transaction with size_i equal to max_val_p uses 0 bits
 *   from the sub-block number since the sub-block is equivalent in size to the whole block.
 *
 *   Consider a system with max_val_p = 7 (8 words per block), where a block comprises words
 *   [7, 6, 5, 4, 3, 2, 1, 0], listed most to least significant. An exampe system like this could
 *   have 512 bit blocks with a stream data width of 64 bits. 3 bits = log2(512/64) are required
 *   for the stream count. The transaction size (size_i) determines how many bits are used from
 *   val_i and cnt_r to produce wrap_o.
 *
 *   E.g., max_val_p = 7 for a system with 512-bit blocks and 64-bit stream data width
 *   A 512-bit transaction sets size_i = 7 and a 256-bit transactions sets size_i = 3
 *   512-bit, size_i = 7, val_i = 2: wrap_o = 2, 3, 4, 5, 6, 7, 0, 1
 *   256-bit, size_i = 3, val_i = 2: wrap_o = 2, 3, 0, 1
 *   512-bit, size_i = 7, val_i = 6: wrap_o = 6, 7, 0, 1, 2, 3, 4, 5
 *   256-bit, size_i = 3, val_i = 6: wrap_o = 6, 7, 4, 5
 *
 */

`include "bsg_defines.v"

module bp_me_wrap_counter
 #(parameter `BSG_INV_PARAM(max_val_p)
   , localparam width_lp = `BSG_WIDTH(max_val_p)
   )
  (input                                          clk_i
   , input                                        reset_i

   // Increment counter
   , input                                        en_i
   // Size of a new transaction
   , input [`BSG_SAFE_MINUS(width_lp,1):0]        size_i
   // Initial value for a new transaction
   , input [`BSG_SAFE_MINUS(width_lp,1):0]        val_i

   // wrap-around count, used to construct proper stream beat address
   // wraps within sub-block aligned portion of block targeted by request
   , output logic [`BSG_SAFE_MINUS(width_lp,1):0] wrap_o
   , output logic                                 first_o
   , output logic                                 last_o
   );

  // parameter check
  if ((max_val_p > 0) && !`BSG_IS_POW2(max_val_p+1))
    $error("max_val_p+1 of %0d is not a power of two...wrap-around counting will break.", max_val_p+1);

  if (max_val_p == 0)
    begin : z
      assign wrap_o = '0;
      assign first_o = 1'b1;
      assign last_o = 1'b1;
    end
  else
    begin : nz
      enum logic {e_ready, e_stream} state_n, state_r;
      wire is_ready = (state_r == e_ready);
      wire is_stream = (state_r == e_stream);
      assign first_o = is_ready;

      logic [width_lp-1:0] cnt_r;
      wire [width_lp-1:0] cnt_val_li = val_i + en_i;
      bsg_counter_set_en
       #(.max_val_p(max_val_p), .reset_val_p('0))
       counter
        (.clk_i(clk_i)
         ,.reset_i(reset_i)

         ,.set_i(is_ready)
         ,.en_i(en_i)
         ,.val_i(cnt_val_li)
         ,.count_o(cnt_r)
         );

      logic [width_lp-1:0] last_cnt_r;
      wire [width_lp-1:0] last_cnt_n = val_i + size_i;
      bsg_dff_en
       #(.width_p(width_lp))
       last_cnt_reg
        (.clk_i(clk_i)
         ,.en_i(is_ready)
         ,.data_i(last_cnt_n)
         ,.data_o(last_cnt_r)
         );
      assign last_o = is_ready ? (size_i == '0) : (last_cnt_r == cnt_r);

      // selection input used to pick bits from block-wrapped and sub-block wrapped counts
      logic [width_lp-1:0] wrap_sel_li;
      for (genvar i = 0; i < width_lp; i++)
        begin : cnt_sel
          assign wrap_sel_li[i] = size_i >= 2**i;
        end

      // sub-block wrapped and aligned count (stream word)
      logic [width_lp-1:0] wrap_lo;
      bsg_mux_bitwise
       #(.width_p(width_lp))
       wrap_mux
        (.data0_i(val_i)
         ,.data1_i(cnt_r)
         ,.sel_i(wrap_sel_li)
         ,.data_o(wrap_lo)
         );

      assign wrap_o = is_ready ? val_i : wrap_lo;

      always_comb begin
        case (state_r)
          e_stream: state_n = (en_i &  last_o) ? e_ready : e_stream;
          // e_ready
          default : state_n = (en_i & ~last_o) ? e_stream : e_ready;
        endcase
      end

      // synopsys sync_set_reset "reset_i"
      always_ff @(posedge clk_i) begin
        if (reset_i) begin
          state_r <= e_ready;
        end else begin
          state_r <= state_n;
        end
      end
    end

endmodule

`BSG_ABSTRACT_MODULE(bp_me_wrap_counter)

