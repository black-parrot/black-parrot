/**
 *
 * Name:
 *   bp_me_cache_slice.sv
 *
 * Description:
 *
 */

`include "bp_common_defines.svh"
`include "bp_me_defines.svh"
`include "bsg_cache.vh"
`include "bsg_noc_links.vh"

module bp_me_cache_slice
 import bp_common_pkg::*;
 import bp_me_pkg::*;
 import bsg_noc_pkg::*;
 import bsg_cache_pkg::*;
 #(parameter bp_params_e bp_params_p = e_bp_default_cfg
   `declare_bp_proc_params(bp_params_p)

   `declare_bp_bedrock_mem_if_widths(paddr_width_p, did_width_p, lce_id_width_p, lce_assoc_p, uce)
   `declare_bp_bedrock_mem_if_widths(paddr_width_p, did_width_p, lce_id_width_p, lce_assoc_p, cce)

   , localparam dma_pkt_width_lp = `bsg_cache_dma_pkt_width(daddr_width_p)
   )
  (input                                                 clk_i
   , input                                               reset_i

   , input  [cce_mem_header_width_lp-1:0]                mem_cmd_header_i
   , input  [l2_data_width_p-1:0]                        mem_cmd_data_i
   , input                                               mem_cmd_v_i
   , output logic                                        mem_cmd_ready_and_o
   , input                                               mem_cmd_last_i

   , output [cce_mem_header_width_lp-1:0]                mem_resp_header_o
   , output [l2_data_width_p-1:0]                        mem_resp_data_o
   , output logic                                        mem_resp_v_o
   , input                                               mem_resp_ready_and_i
   , output logic                                        mem_resp_last_o

   // DRAM interface
   , output logic [l2_banks_p-1:0][dma_pkt_width_lp-1:0] dma_pkt_o
   , output logic [l2_banks_p-1:0]                       dma_pkt_v_o
   , input [l2_banks_p-1:0]                              dma_pkt_ready_and_i

   , input [l2_banks_p-1:0][l2_fill_width_p-1:0]         dma_data_i
   , input [l2_banks_p-1:0]                              dma_data_v_i
   , output logic [l2_banks_p-1:0]                       dma_data_ready_and_o

   , output logic [l2_banks_p-1:0][l2_fill_width_p-1:0]  dma_data_o
   , output logic [l2_banks_p-1:0]                       dma_data_v_o
   , input [l2_banks_p-1:0]                              dma_data_ready_and_i
   );

  `declare_bp_cfg_bus_s(hio_width_p, core_id_width_p, cce_id_width_p, lce_id_width_p);
  `declare_bp_bedrock_mem_if(paddr_width_p, did_width_p, lce_id_width_p, lce_assoc_p, uce);

  `declare_bsg_cache_pkt_s(daddr_width_p, l2_data_width_p);
  bsg_cache_pkt_s [l2_banks_p-1:0] cache_pkt_li;
  logic [l2_banks_p-1:0] cache_pkt_v_li, cache_pkt_ready_and_lo;
  logic [l2_banks_p-1:0][l2_data_width_p-1:0] cache_data_lo;
  logic [l2_banks_p-1:0] cache_data_v_lo, cache_data_ready_and_li;

  bp_me_cce_to_cache
   #(.bp_params_p(bp_params_p))
   cce_to_cache
    (.clk_i(clk_i)
     ,.reset_i(reset_i)

     ,.mem_cmd_header_i(mem_cmd_header_i)
     ,.mem_cmd_data_i(mem_cmd_data_i)
     ,.mem_cmd_v_i(mem_cmd_v_i)
     ,.mem_cmd_ready_and_o(mem_cmd_ready_and_o)
     ,.mem_cmd_last_i(mem_cmd_last_i)

     ,.mem_resp_header_o(mem_resp_header_o)
     ,.mem_resp_data_o(mem_resp_data_o)
     ,.mem_resp_v_o(mem_resp_v_o)
     ,.mem_resp_ready_and_i(mem_resp_ready_and_i)
     ,.mem_resp_last_o(mem_resp_last_o)

     ,.cache_pkt_o(cache_pkt_li)
     ,.cache_pkt_v_o(cache_pkt_v_li)
     ,.cache_pkt_ready_and_i(cache_pkt_ready_and_lo)

     ,.cache_data_i(cache_data_lo)
     ,.cache_data_v_i(cache_data_v_lo)
     ,.cache_data_yumi_o(cache_data_yumi_li)
     );

  for (genvar i = 0; i < l2_banks_p; i++)
    begin : bank
      bsg_cache
       #(.addr_width_p(daddr_width_p)
         ,.data_width_p(l2_data_width_p)
         ,.dma_data_width_p(l2_fill_width_p)
         ,.block_size_in_words_p(l2_block_size_in_words_p)
         ,.sets_p((l2_banks_p > 0) ? l2_sets_p : 2)
         ,.ways_p((l2_banks_p > 0) ? l2_assoc_p : 2)
         ,.amo_support_p(((l2_amo_support_p[e_amo_swap]) << e_cache_amo_swap)
                         | ((l2_amo_support_p[e_amo_fetch_logic]) << e_cache_amo_xor)
                         | ((l2_amo_support_p[e_amo_fetch_logic]) << e_cache_amo_and)
                         | ((l2_amo_support_p[e_amo_fetch_logic]) << e_cache_amo_or)
                         | ((l2_amo_support_p[e_amo_fetch_arithmetic]) << e_cache_amo_add)
                         | ((l2_amo_support_p[e_amo_fetch_arithmetic]) << e_cache_amo_min)
                         | ((l2_amo_support_p[e_amo_fetch_arithmetic]) << e_cache_amo_max)
                         | ((l2_amo_support_p[e_amo_fetch_arithmetic]) << e_cache_amo_minu)
                         | ((l2_amo_support_p[e_amo_fetch_arithmetic]) << e_cache_amo_maxu)
                         )
        )
       cache
        (.clk_i(clk_i)
         ,.reset_i(reset_i)

         ,.cache_pkt_i(cache_pkt_li[i])
         ,.v_i(cache_pkt_v_li[i])
         ,.ready_o(cache_pkt_ready_and_lo[i])

         ,.data_o(cache_data_lo[i])
         ,.v_o(cache_data_v_lo[i])
         ,.yumi_i(cache_data_yumi_li[i])

         ,.dma_pkt_o(dma_pkt_o[i])
         ,.dma_pkt_v_o(dma_pkt_v_o[i])
         ,.dma_pkt_yumi_i(dma_pkt_ready_and_i[i] & dma_pkt_v_o[i])

         ,.dma_data_i(dma_data_i[i])
         ,.dma_data_v_i(dma_data_v_i[i])
         ,.dma_data_ready_o(dma_data_ready_and_o[i])

         ,.dma_data_o(dma_data_o[i])
         ,.dma_data_v_o(dma_data_v_o[i])
         ,.dma_data_yumi_i(dma_data_ready_and_i[i] & dma_data_v_o[i])

         ,.v_we_o()
         );
    end

  // TODO: Wrap
  logic l2_clk_lo, l2_reset_lo;
  localparam l2_ds_width_lp = `BSG_WIDTH(l2_downclock_p/2);
  if (l2_downclock_p > 1)
    begin : dc
      bsg_counter_clock_downsample
       #(.width_p(l2_ds_width_lp))
       l2_ds
        (.clk_i(clk_i)
         ,.reset_i(reset_i)

         ,.val_i(l2_ds_width_lp'(l2_downclock_p/2-1))
         ,.clk_r_o(l2_clk_lo)
         );

      bsg_dff_chain
       #(.width_p(1), .num_stages_p(2*l2_downclock_p-1))
       l2_reset_chain
        (.clk_i(clk_i)
         ,.data_i(reset_i)
         ,.data_o(l2_reset_lo)
         );
    end
  else
    begin : ndc
      assign l2_clk_lo = clk_i;
      assign l2_reset_lo = reset_i;
    end

  logic l2_pkt_v_li, l2_pkt_ready_lo;
  logic l2_dma_data_v_li, l2_dma_data_ready_lo;
  bsg_fifo_1r1w_periodic
   #(.a_period_p(1), .b_period_p(l2_downclock_p), .num_hs_p(2))
   cache_downclock
    (.a_clk_i(clk_i)
     ,.a_reset_i(reset_i)
     ,.a_v_i({cache_pkt_v_li, dma_data_v_i})
     ,.a_ready_and_o({cache_pkt_ready_and_lo, dma_data_ready_and_o})

     ,.b_clk_i(l2_clk_lo)
     ,.b_reset_i(l2_reset_lo)
     ,.b_v_o({l2_pkt_v_li, l2_dma_data_v_li})
     ,.b_ready_and_i({l2_pkt_ready_lo, l2_dma_data_ready_lo})
     );

  logic l2_data_v_lo, l2_data_ready_and_li;
  logic l2_dma_pkt_v_lo, l2_dma_pkt_ready_and_li;
  logic l2_dma_data_v_lo, l2_dma_data_ready_and_li;
  bsg_fifo_1r1w_periodic
   #(.a_period_p(l2_downclock_p), .b_period_p(1), .num_hs_p(3))
   cache_upclock
    (.a_clk_i(l2_clk_lo)
     ,.a_reset_i(l2_reset_lo)
     ,.a_v_i({l2_data_v_lo, l2_dma_pkt_v_lo, l2_dma_data_v_lo})
     ,.a_ready_and_o({l2_data_ready_and_li, l2_dma_pkt_ready_and_li, l2_dma_data_ready_and_li})

     ,.b_clk_i(clk_i)
     ,.b_reset_i(reset_i)
     ,.b_v_o({cache_data_v_lo, dma_pkt_v_o, dma_data_v_o})
     ,.b_ready_and_i({cache_data_ready_and_li, dma_pkt_yumi_i, dma_data_yumi_i})
     );

endmodule

