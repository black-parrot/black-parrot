package pc_gen_pkg;


endpackage : pc_gen_pkg
