
package bp_fe_pkg;

endpackage

