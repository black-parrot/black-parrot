
package bp_top_pkg;

endpackage

