/**
 *  Name:
 *    bp_be_dcache_pkg.vh
 *  
 *  Description:
 *    opcodes for dcache packet from mmu.
 */

package bp_be_dcache_pkg;
    
  `include "bp_be_dcache_pkt.vh"
  `include "bp_be_dcache_pipeline.vh"
  `include "bp_be_dcache_tag_info.vh"
  `include "bp_be_dcache_wbuf_entry.vh"
  `include "../bp_be_ctl_defines.vh"

endpackage
