/*
 * bp_me_pkg.svh
 *
 * Contains the interface structures used for communicating between the CCE and Memory.
 *
 */

package bp_me_pkg;

  import bp_common_pkg::*;

  `include "bp_me_cce_pkgdef.svh"
  `include "bp_me_cce_inst_pkgdef.svh"
  `include "bp_me_axi_pkgdef.sv"

endpackage

