
`ifndef BP_COMMON_CACHE_PKGDEF_SVH
`define BP_COMMON_CACHE_PKGDEF_SVH

  localparam cache_base_addr_gp        = 'h0400_0000;
  localparam cache_tagfl_base_addr_gp  = 20'h0_0000;

`endif

