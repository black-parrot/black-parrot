/**
 *  Name:
 *    bp_be_dcache_pkg.svh
 *
 *  Description:
 *    opcodes for dcache packet from mmu.
 */

package bp_be_dcache_pkg;

  `include "bp_be_dcache_pkt.svh"
  `include "bp_be_dcache_pipeline.svh"
  `include "bp_be_dcache_tag_info.svh"
  `include "bp_be_dcache_wbuf_entry.svh"
  `include "bp_be_ctl_defines.svh"

endpackage
