`ifndef BP_ME_DEFINES_SVH
`define BP_ME_DEFINES_SVH

  `include "bp_me_cache_defines.svh"
  `include "bp_me_cce_defines.svh"
  `include "bp_me_cce_inst_defines.svh"
  `include "bp_me_wormhole_defines.svh"

`endif

