
package bp_fe_pkg;

  `include "bsg_defines.v"
  `include "bp_common_core_if.vh"
  `include "bp_fe_defines.vh"
  `include "bp_fe_mem_defines.vh"

endpackage : bp_fe_pkg
