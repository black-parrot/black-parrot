
`ifndef BP_COMMON_CLINT_PKGDEF_SVH
`define BP_COMMON_CLINT_PKGDEF_SVH

  localparam clint_base_addr_gp        = 'h0300_0000;
  localparam mipi_reg_base_addr_gp     = 32'h0030_0000;
  localparam mtimecmp_reg_base_addr_gp = 32'h0030_4000;
  localparam mtime_reg_addr_gp         = 32'h0030_bff8;
  localparam plic_reg_base_addr_gp     = 32'h0030_b000;

`endif

