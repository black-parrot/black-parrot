
package bp_fe_pkg;

  `include "bp_fe_icache_pkgdef.svh"
  `include "bp_fe_pc_gen_pkgdef.svh"

endpackage

