/**
 * bp_me_nonsynth_mock_lce.v
 *
 * This mock LCE behaves like a mock D$. It connects to a trace replay module and to the BP ME.
 * The trace replay format is the same as the trace replay format for the D$.
 */

module tag_lookup
  import bp_common_pkg::*;
  #(parameter lce_assoc_p="inv"
    , parameter ptag_width_p="inv"
    , parameter coh_bits_p="inv"
    , localparam tag_s_width_lp=(coh_bits_p+ptag_width_p)
    , localparam lg_lce_assoc_lp=`BSG_SAFE_CLOG2(lce_assoc_p)
   )
  (input [lce_assoc_p-1:0][tag_s_width_lp-1:0] tag_set_i
   , input [ptag_width_p-1:0] ptag_i
   , output logic hit_o
   , output logic dirty_o
   , output logic [lg_lce_assoc_lp-1:0] way_o
   , input [lg_lce_assoc_lp-1:0] lru_way_i
   , output logic lru_dirty_o
  );
  typedef struct packed {
    logic [coh_bits_p-1:0] coh_st;
    logic [ptag_width_p-1:0] tag;
  } tag_s;

  tag_s [lce_assoc_p-1:0] tags;
  assign tags = tag_set_i;

  logic [lce_assoc_p-1:0] hits;
  int i;
  always_comb begin
    for (i = 0; i < lce_assoc_p; i=i+1) begin
      if (tags[i].tag == ptag_i && tags[i].coh_st != e_MESI_I) begin
        hits[i] = 1'b1;
      end else begin
        hits[i] = '0;
      end
    end
  end

  bsg_encode_one_hot
    #(.width_p(lce_assoc_p))
  hits_to_way_id
    (.i(hits)
     ,.addr_o(way_o)
     ,.v_o(hit_o)
    );

  assign dirty_o = (tags[way_o].coh_st == e_MESI_M);
  assign lru_dirty_o = (tags[lru_way_i].coh_st == e_MESI_M);

endmodule


module bp_me_nonsynth_mock_lce
  import bp_common_pkg::*;
  import bp_common_aviary_pkg::*;
  import bp_cce_pkg::*;
  import bp_be_dcache_pkg::*;
  #(parameter bp_cfg_e cfg_p = e_bp_half_core_cfg
    `declare_bp_proc_params(cfg_p)

    , localparam block_size_in_bytes_lp=(cce_block_width_p / 8)

    , localparam dcache_opcode_width_lp=$bits(bp_be_dcache_opcode_e)
    , localparam tr_ring_width_lp=(dcache_opcode_width_lp+paddr_width_p+dword_width_p)

    , localparam block_offset_bits_lp=`BSG_SAFE_CLOG2(block_size_in_bytes_lp)

    , localparam lg_lce_sets_lp=`BSG_SAFE_CLOG2(lce_sets_p)
    , localparam lg_lce_assoc_lp=`BSG_SAFE_CLOG2(lce_assoc_p)
    , localparam lg_num_lce_lp=`BSG_SAFE_CLOG2(num_lce_p)
    , localparam lg_num_cce_lp=`BSG_SAFE_CLOG2(num_cce_p)

    , localparam ptag_width_lp=paddr_width_p-lg_lce_sets_lp-block_offset_bits_lp

`declare_bp_lce_cce_if_widths(num_cce_p, num_lce_p, paddr_width_p, lce_assoc_p, dword_width_p, cce_block_width_p)
  )
  (
    input                                                   clk_i
    ,input                                                  reset_i

    ,input [lg_num_lce_lp-1:0]                              lce_id_i

    // the input packets are the same as the dcache trace replay packets: {dcache_cmd, paddr, data}
    ,input [tr_ring_width_lp-1:0]                           tr_pkt_i
    ,input                                                  tr_pkt_v_i
    ,output logic                                           tr_pkt_yumi_o

    ,output logic [tr_ring_width_lp-1:0]                    tr_pkt_o
    ,output logic                                           tr_pkt_v_o
    ,input                                                  tr_pkt_ready_i

    // LCE-CCE Interface
    // inbound: valid->ready (a.k.a. valid->yumi), demanding
    // outbound: ready->valid, demanding
    ,output logic [lce_cce_req_width_lp-1:0]                lce_req_o
    ,output logic                                           lce_req_v_o
    ,input                                                  lce_req_ready_i

    ,output logic [lce_cce_resp_width_lp-1:0]               lce_resp_o
    ,output logic                                           lce_resp_v_o
    ,input                                                  lce_resp_ready_i

    ,output logic [lce_cce_data_resp_width_lp-1:0]          lce_data_resp_o
    ,output logic                                           lce_data_resp_v_o
    ,input                                                  lce_data_resp_ready_i

    ,input [cce_lce_cmd_width_lp-1:0]                       lce_cmd_i
    ,input                                                  lce_cmd_v_i
    ,output logic                                           lce_cmd_ready_o

    ,input [lce_data_cmd_width_lp-1:0]                      lce_data_cmd_i
    ,input                                                  lce_data_cmd_v_i
    ,output logic                                           lce_data_cmd_ready_o

    ,output logic [lce_data_cmd_width_lp-1:0]               lce_data_cmd_o
    ,output logic                                           lce_data_cmd_v_o
    ,input                                                  lce_data_cmd_ready_i
  );

  // LCE-CCE interface structs
  `declare_bp_lce_cce_if(num_cce_p, num_lce_p, paddr_width_p, lce_assoc_p, dword_width_p, cce_block_width_p);

  // Structs for output messages
  bp_lce_cce_req_s lce_req_s;
  bp_lce_cce_resp_s lce_resp_s;
  bp_lce_cce_data_resp_s lce_data_resp_s;
  bp_lce_data_cmd_s lce_data_cmd_s;
  assign lce_req_o = lce_req_s;
  assign lce_resp_o = lce_resp_s;
  assign lce_data_resp_o = lce_data_resp_s;
  assign lce_data_cmd_o = lce_data_cmd_s;

  // FIFO to buffer LCE commands from ME
  logic lce_cmd_v, lce_cmd_yumi;
  logic [cce_lce_cmd_width_lp-1:0] lce_cmd_bits;
  bp_cce_lce_cmd_s lce_cmd, lce_cmd_r, lce_cmd_n;
  assign lce_cmd = lce_cmd_bits;

  bsg_two_fifo
    #(.width_p(cce_lce_cmd_width_lp))
  lce_cmd_fifo
    (.clk_i(clk_i)
     ,.reset_i(reset_i)
     // to/from ME
     ,.ready_o(lce_cmd_ready_o)
     ,.data_i(lce_cmd_i)
     ,.v_i(lce_cmd_v_i)
     // to/from mock LCE
     ,.v_o(lce_cmd_v)
     ,.data_o(lce_cmd_bits)
     ,.yumi_i(lce_cmd_yumi)
    );

  // FIFO to buffer LCE Data commands from ME
  logic lce_data_cmd_v, lce_data_cmd_yumi;
  logic [lce_data_cmd_width_lp-1:0] lce_data_cmd_bits;
  bp_lce_data_cmd_s lce_data_cmd, lce_data_cmd_r, lce_data_cmd_n;
  assign lce_data_cmd = lce_data_cmd_bits;

  bsg_two_fifo
    #(.width_p(lce_data_cmd_width_lp))
  lce_data_cmd_fifo
    (.clk_i(clk_i)
     ,.reset_i(reset_i)
     // to/from ME
     ,.ready_o(lce_data_cmd_ready_o)
     ,.data_i(lce_data_cmd_i)
     ,.v_i(lce_data_cmd_v_i)
     // to/from mock LCE
     ,.v_o(lce_data_cmd_v)
     ,.data_o(lce_data_cmd_bits)
     ,.yumi_i(lce_data_cmd_yumi)
    );

////////////////////////////////////////////////////////////////////////////////////////////////////
// Tag and Data arrays
////////////////////////////////////////////////////////////////////////////////////////////////////

  typedef struct packed {
    logic [`bp_cce_coh_bits-1:0] coh_st;
    logic [ptag_width_lp-1:0] tag;
  } tag_s;

  localparam tag_s_width_lp = $bits(tag_s);

  // Tags
  tag_s [lce_sets_p-1:0][lce_assoc_p-1:0] tags, tag_n;
  logic [lce_sets_p-1:0][lce_assoc_p-1:0] tag_w;
  always_ff @(posedge clk_i) begin
    for (integer i = 0; i < lce_sets_p; i=i+1) begin
      for (integer j = 0; j < lce_assoc_p; j=j+1) begin
        if (tag_w[i][j]) begin
          tags[i][j] <= tag_n[i][j];
        end
      end
    end
  end

  // async read of tags at specified set and way
  tag_s tag_cur;
  logic [lg_lce_sets_lp-1:0] tag_set;
  logic [lg_lce_assoc_lp-1:0] tag_way;
  assign tag_cur = tags[tag_set][tag_way];

  // Data
  logic [lce_sets_p-1:0][lce_assoc_p-1:0][cce_block_width_p-1:0] data, data_n, data_mask_n;
  logic [lce_sets_p-1:0][lce_assoc_p-1:0] data_w;
  always_ff @(posedge clk_i) begin
    for (integer i = 0; i < lce_sets_p; i=i+1) begin
      for (integer j = 0; j < lce_assoc_p; j=j+1) begin
        if (data_w[i][j]) begin
          for (integer k = 0; k < cce_block_width_p; k=k+1) begin
            if (data_mask_n[k]) begin
              data[i][j][k] <= data_n[k];
            end
          end
        end
      end
    end
  end

  // async read of data at specified set and way
  logic [cce_block_width_p-1:0] data_cur;
  logic [lg_lce_sets_lp-1:0] data_set;
  logic [lg_lce_assoc_lp-1:0] data_way;
  assign data_cur = data[data_set][data_way];


////////////////////////////////////////////////////////////////////////////////////////////////////
// Trace Replay Command
////////////////////////////////////////////////////////////////////////////////////////////////////

  // current command from trace replay
  typedef struct packed {
    logic [dcache_opcode_width_lp-1:0] cmd;
    logic [paddr_width_p-1:0]          paddr;
    logic [dword_width_p-1:0]          data;
  } tr_cmd_s;

  // current command being processed
  tr_cmd_s cmd, cmd_n;
  always_ff @(posedge clk_i) begin
    if (reset_i) begin
      cmd <= '0;
    end else begin
      cmd <= cmd_n;
    end
  end

  // some useful signals from the current trace replay command
  logic store_op, load_op, signed_op, byte_op, word_op, double_op, half_op;
  logic [1:0] op_size;
  logic [2:0] dword_offset;
  logic [2:0] byte_offset;
  assign store_op = cmd.cmd[3];
  assign load_op = ~cmd.cmd[3];
  assign signed_op = ~cmd.cmd[2];
  assign op_size = cmd.cmd[1:0];
  assign double_op = (cmd.cmd[1:0] == 2'b11);
  assign word_op = (cmd.cmd[1:0] == 2'b10);
  assign half_op = (cmd.cmd[1:0] == 2'b01);
  assign byte_op = (cmd.cmd[1:0] == 2'b00);
  assign dword_offset = cmd.paddr[5:3];
  assign byte_offset = cmd.paddr[2:0];

  // Data word (64-bit) targeted by current trace replay command
  logic [dword_width_p-1:0] load_data;
  assign load_data = data_cur[dword_width_p*dword_offset +: dword_width_p];
  logic word_sigext, half_sigext, byte_sigext;
  logic [31:0] load_word;
  logic [15:0] load_half;
  logic [7:0] load_byte;

  bsg_mux #(
    .width_p(32)
    ,.els_p(2)
  ) word_mux (
    .data_i(load_data)
    ,.sel_i(byte_offset[2])
    ,.data_o(load_word)
  );
  
  bsg_mux #(
    .width_p(16)
    ,.els_p(4)
  ) half_mux (
    .data_i(load_data)
    ,.sel_i(byte_offset[2:1])
    ,.data_o(load_half)
  );

  bsg_mux #(
    .width_p(8)
    ,.els_p(8)
  ) byte_mux (
    .data_i(load_data)
    ,.sel_i(byte_offset[2:0])
    ,.data_o(load_byte)
  );

  assign word_sigext = signed_op & load_word[31]; 
  assign half_sigext = signed_op & load_half[15]; 
  assign byte_sigext = signed_op & load_byte[7]; 

  // Tag lookup
  // inputs
  tag_s [lce_assoc_p-1:0] tag_set_li;
  logic [ptag_width_lp-1:0] ptag_li;
  logic [lg_lce_assoc_lp-1:0] lru_way_r, lru_way_n, lru_way_li;
  // outputs
  logic tag_hit_r, tag_hit_n, tag_hit_lo;
  logic tag_dirty_r, tag_dirty_n, tag_dirty_lo;
  logic [lg_lce_assoc_lp-1:0] tag_hit_way_r, tag_hit_way_n, tag_hit_way_lo;
  logic lru_dirty_r, lru_dirty_n, lru_dirty_lo;

  always_ff @(posedge clk_i) begin
    if (reset_i) begin
      lru_way_r <= '0;
      tag_hit_r <= '0;
      tag_dirty_r <= '0;
      tag_hit_way_r <= '0;
      lru_dirty_r <= '0;
    end else begin
      lru_way_r <= lru_way_n;
      tag_hit_r <= tag_hit_n;
      tag_dirty_r <= tag_dirty_n;
      tag_hit_way_r <= tag_hit_way_n;
      lru_dirty_r <= lru_dirty_n;
    end
  end

  tag_lookup
    #(.lce_assoc_p(lce_assoc_p)
      ,.ptag_width_p(ptag_width_lp)
      ,.coh_bits_p(`bp_cce_coh_bits)
      )
  lce_tag_lookup
    (.tag_set_i(tag_set_li)
     ,.ptag_i(ptag_li)
     ,.lru_way_i(lru_way_li)
     ,.hit_o(tag_hit_lo)
     ,.dirty_o(tag_dirty_lo)
     ,.way_o(tag_hit_way_lo)
     ,.lru_dirty_o(lru_dirty_lo)
     );

  typedef enum logic [7:0] {
    RESET
    ,SET_CLEAR
    ,SYNC
    ,READY

    ,LCE_DATA_CMD
    ,LCE_DATA_CMD_WR_DATA

    ,LCE_CMD
    ,LCE_CMD_TR
    ,LCE_CMD_WB
    ,LCE_CMD_INV
    ,LCE_CMD_INV_RESP
    ,LCE_CMD_ST
    ,LCE_CMD_STW
    ,LCE_CMD_STW_RESP

    ,LCE_CMD_ST_DATA_RESP

    ,TR_CMD
    ,TR_CMD_LD_HIT
    ,TR_CMD_LD_MISS
    ,TR_CMD_ST_HIT
    ,TR_CMD_ST_HIT_RESP
    ,TR_CMD_ST_MISS

    ,FINISH_MISS
  } lce_state_e;

  lce_state_e lce_state, lce_state_n;

  // miss handling state
  logic miss_r, miss_n;
  logic [lg_lce_assoc_lp-1:0] miss_lru_way_r, miss_lru_way_n;
  logic miss_st_upgrade_r, miss_st_upgrade_n;
  logic tag_received_r, tag_received_n;
  logic data_received_r, data_received_n;

  always_ff @(posedge clk_i) begin
    if (reset_i) begin
      lce_state <= RESET;

      lce_cmd_r <= '0;
      lce_data_cmd_r <= '0;

      miss_r <= '0;
      miss_lru_way_r <= '0;
      miss_st_upgrade_r <= '0;
      tag_received_r <= '0;
      data_received_r <= '0;

    end else begin
      lce_state <= lce_state_n;

      lce_cmd_r <= lce_cmd_n;
      lce_data_cmd_r <= lce_data_cmd_n;

      miss_r <= miss_n;
      miss_lru_way_r <= miss_lru_way_n;
      miss_st_upgrade_r <= miss_st_upgrade_n;
      tag_received_r <= tag_received_n;
      data_received_r <= data_received_n;

    end
  end


  always_comb begin
    if (reset_i) begin
      lce_state_n = RESET;

      // trace replay command inbound
      cmd_n = '0;
      tr_pkt_yumi_o = '0;

      // trace replay response out
      tr_pkt_o = '0;
      tr_pkt_v_o = '0;

      // outbound queues
      lce_req_v_o = '0;
      lce_req_s = '0;
      lce_resp_v_o = '0;
      lce_resp_s = '0;
      lce_data_resp_v_o = '0;
      lce_data_resp_s = '0;
      lce_data_cmd_v_o = '0;
      lce_data_cmd_s = '0;

      // inbound queues
      lce_cmd_n = '0;
      lce_cmd_yumi = '0;
      lce_data_cmd_n ='0;
      lce_data_cmd_yumi = '0;

      // miss handling
      lru_way_n = '0;
      miss_n = '0;
      miss_lru_way_n = '0;
      miss_st_upgrade_n = '0;
      tag_received_n = '0;
      data_received_n = '0;

      // tag and data arrays
      tag_n = '0;
      tag_w = '0;
      data_n = '0;
      data_w = '0;
      data_mask_n = '0;

      // tag lookup module
      tag_set_li = '0;
      ptag_li = '0;
      lru_way_li = '0;
      lru_way_n = '0;
      tag_hit_n = '0;
      tag_dirty_n = '0;
      tag_hit_way_n = '0;
      lru_dirty_n = '0;

      // other stuff
      tag_set = '0;
      tag_way = '0;
      data_set = '0;
      data_way = '0;

    end else begin
      lce_state_n = RESET;

      // trace replay command inbound
      cmd_n = cmd;
      tr_pkt_yumi_o = '0;

      // trace replay response out
      tr_pkt_o = '0;
      tr_pkt_v_o = '0;

      // outbound queues
      lce_req_v_o = '0;
      lce_req_s = '0;
      lce_resp_v_o = '0;
      lce_resp_s = '0;
      lce_data_resp_v_o = '0;
      lce_data_resp_s = '0;
      lce_data_cmd_v_o = '0;
      lce_data_cmd_s = '0;

      // inbound queues
      lce_cmd_n = lce_cmd_r;
      lce_cmd_yumi = '0;
      lce_data_cmd_n =lce_data_cmd_r;
      lce_data_cmd_yumi = '0;

      // miss handling
      lru_way_n = lru_way_r;
      miss_n = miss_r;
      miss_lru_way_n = miss_lru_way_r;
      miss_st_upgrade_n = miss_st_upgrade_r;
      tag_received_n = tag_received_r;
      data_received_n = data_received_r;

      // tag and data arrays
      tag_n = '0;
      tag_w = '0;
      data_n = '0;
      data_w = '0;
      data_mask_n = '0;

      // tag lookup module
      tag_set_li = '0;
      ptag_li = '0;
      lru_way_li = '0;
      lru_way_n = lru_way_r;
      tag_hit_n = tag_hit_r;
      tag_dirty_n = tag_dirty_r;
      tag_hit_way_n = tag_hit_way_r;
      lru_dirty_n = lru_dirty_r;

      // other stuff
      tag_set = '0;
      tag_way = '0;
      data_set = '0;
      data_way = '0;

      case (lce_state)
        RESET: begin
          lce_state_n = SET_CLEAR;
        end
        SET_CLEAR: begin
          // by default, stay in SET_CLEAR, waiting for set clear commands to arrive
          lce_state_n = SET_CLEAR;

          if (lce_cmd_v && lce_cmd.msg_type == e_lce_cmd_sync) begin
            // dequeue the command, go to SYNC
            lce_cmd_yumi = 1'b1;
            lce_cmd_n = lce_cmd;
            lce_state_n = SYNC;
          end else if (lce_cmd_v && lce_cmd.msg_type == e_lce_cmd_set_clear) begin
            // dequeue the command
            lce_cmd_yumi = 1'b1;
            lce_cmd_n = lce_cmd;

            // clear set in cache
            tag_w[tag_set] = '1;
            tag_n[tag_set] = '0;

            lce_state_n = SET_CLEAR;
          end
        end
        SYNC: begin
          // create the LCE response and make it valid for output
          lce_resp_s.dst_id = lce_cmd_r.src_id;
          lce_resp_s.src_id = lce_id_i;
          lce_resp_s.msg_type = e_lce_cce_sync_ack;
          lce_resp_s.addr = '0;
          lce_resp_v_o = 1'b1;

          // response goes out if inbound ready signal is high (ready&valid)
          lce_state_n = (lce_resp_ready_i) ? READY : SYNC;
        end
        READY: begin
          lce_state_n = READY;
          if (lce_data_cmd_v) begin
            lce_data_cmd_yumi = 1'b1;
            lce_data_cmd_n = lce_data_cmd;
            lce_state_n = LCE_DATA_CMD;
          end else if (lce_cmd_v) begin
            // dequeue the command and save
            lce_cmd_yumi = 1'b1;
            lce_cmd_n = lce_cmd;
            if (lce_cmd.msg_type == e_lce_cmd_invalidate_tag) begin
              lce_state_n = LCE_CMD_INV;
            end else if (lce_cmd.msg_type == e_lce_cmd_transfer) begin
              lce_state_n = LCE_CMD_TR;
            end else if (lce_cmd.msg_type == e_lce_cmd_writeback) begin
              lce_state_n = LCE_CMD_WB;
            end else if (lce_cmd.msg_type == e_lce_cmd_set_tag) begin
              lce_state_n = LCE_CMD_ST;
            end else if (lce_cmd.msg_type == e_lce_cmd_set_tag_wakeup) begin
              lce_state_n = LCE_CMD_STW;
            end else begin
              lce_state_n = RESET;
              $error("unrecognized LCE command received");
            end

          end else if (tr_pkt_v_i & ~miss_r) begin
            // only process a new trace replay request if not already missing
            tr_pkt_yumi_o = 1'b1;
            cmd_n = tr_pkt_i;
            lce_state_n = TR_CMD;
          end

        end
        LCE_DATA_CMD: begin
          // write the full cache block to data array
          data_mask_n = '1;
          data_set = cmd.paddr[block_offset_bits_lp +: lg_lce_sets_lp];
          data_way = lce_data_cmd_r.way_id;
          data_w[data_set][data_way] = '1;
          data_n = lce_data_cmd.data;
          data_received_n = 1'b1;

          // if tag already received, next state will send response, otherwise wait for tag
          lce_state_n = (tag_received_r) ? LCE_CMD_ST_DATA_RESP : READY;
        end
        LCE_CMD_INV: begin
          // invalidate cmd received - update tags
          tag_set = lce_cmd_r.addr[block_offset_bits_lp +: lg_lce_sets_lp];
          tag_way = lce_cmd_r.way_id;
          tag_w[tag_set][tag_way] = 1'b1;
          tag_n[tag_set][tag_way].coh_st = e_MESI_I;
          tag_n[tag_set][tag_way].tag = lce_cmd_r.addr[paddr_width_p-1 -: ptag_width_lp];

          // send inv_ack next
          lce_state_n = LCE_CMD_INV_RESP;

        end
        LCE_CMD_INV_RESP: begin
          // make the LCE response valid
          lce_resp_s.dst_id = lce_cmd_r.src_id;
          lce_resp_s.src_id = lce_id_i;
          lce_resp_s.msg_type = e_lce_cce_inv_ack;
          lce_resp_s.addr = lce_cmd_r.addr;
          lce_resp_v_o = 1'b1;

          // wait until response accepted (r&v) then go to READY
          lce_state_n = (lce_resp_ready_i) ? READY : LCE_CMD_INV_RESP;

        end
        LCE_CMD_TR: begin
          // transfer cmd

          // data select
          data_set = lce_cmd_r.addr[block_offset_bits_lp +: lg_lce_sets_lp];
          data_way = lce_cmd_r.way_id;

          lce_data_cmd_s.data = data_cur;
          lce_data_cmd_s.dst_id = lce_cmd_r.target;
          lce_data_cmd_s.msg_type = e_lce_data_cmd_transfer;
          lce_data_cmd_s.way_id = lce_cmd_r.target_way_id;
          lce_data_cmd_v_o = 1'b1;

          // wait until data commmand out accepted (r&v), then go to ready
          lce_state_n = (lce_data_cmd_ready_i) ? READY : LCE_CMD_TR;

        end
        LCE_CMD_WB: begin
          // writeback cmd

          // tag and data select
          tag_set = lce_cmd_r.addr[block_offset_bits_lp +: lg_lce_sets_lp];
          tag_way = lce_cmd_r.way_id;
          data_set = lce_cmd_r.addr[block_offset_bits_lp +: lg_lce_sets_lp];
          data_way = lce_cmd_r.way_id;

          if (tag_cur.coh_st == e_MESI_M) begin
            lce_data_resp_s.data = data_cur;
            lce_data_resp_s.msg_type = e_lce_resp_wb;
          end else begin
            lce_data_resp_s.data = '0;
            lce_data_resp_s.msg_type = e_lce_resp_null_wb;
          end
          lce_data_resp_s.dst_id = lce_cmd_r.src_id;
          lce_data_resp_s.src_id = lce_id_i;
          lce_data_resp_s.addr = lce_cmd_r.addr;
          lce_data_resp_v_o = 1'b1;

          // wait until data response accepted (r&v), then go to ready
          lce_state_n = (lce_data_resp_ready_i) ? READY : LCE_CMD_WB;

        end
        LCE_CMD_ST: begin
          // response to miss - tag
          tag_set = lce_cmd_r.addr[block_offset_bits_lp +: lg_lce_sets_lp];
          tag_way = lce_cmd_r.way_id;
          tag_w[tag_set][tag_way] = 1'b1;
          tag_n[tag_set][tag_way].coh_st = lce_cmd_r.state;
          tag_n[tag_set][tag_way].tag = lce_cmd_r.addr[paddr_width_p-1 -: ptag_width_lp];

          tag_received_n = 1'b1;

          // if data already received, send coh_ack or tr_ack next, else wait for data
          lce_state_n = (data_received_r) ? LCE_CMD_ST_DATA_RESP : READY;

        end
        LCE_CMD_ST_DATA_RESP: begin
          lce_resp_s.dst_id = lce_cmd_r.src_id;
          lce_resp_s.src_id = lce_id_i;
          lce_resp_s.msg_type = (lce_data_cmd_r.msg_type == e_lce_data_cmd_transfer) ? e_lce_cce_tr_ack : e_lce_cce_coh_ack;
          lce_resp_s.addr = lce_cmd_r.addr;
          lce_resp_v_o = 1'b1;

          // send ack in response to tag and data both received
          // then, send response back to trace replay
          lce_state_n = (lce_resp_ready_i) ? FINISH_MISS : LCE_CMD_ST_DATA_RESP;
        end
        LCE_CMD_STW: begin
          // update tag array
          tag_set = lce_cmd_r.addr[block_offset_bits_lp +: lg_lce_sets_lp];
          tag_way = lce_cmd_r.way_id;
          tag_w[tag_set][tag_way] = 1'b1;
          tag_n[tag_set][tag_way].coh_st = lce_cmd_r.state;
          tag_n[tag_set][tag_way].tag = lce_cmd_r.addr[paddr_width_p-1 -: ptag_width_lp];

          // send coh_ack next cycle
          lce_state_n = LCE_CMD_STW_RESP;

        end
        LCE_CMD_STW_RESP: begin
          // Send coherence ack in response to set tag and wakeup
          lce_resp_s.dst_id = lce_cmd_r.src_id;
          lce_resp_s.src_id = lce_id_i;
          lce_resp_s.msg_type = e_lce_cce_coh_ack;
          lce_resp_s.addr = lce_cmd_r.addr;
          lce_resp_v_o = 1'b1;

          // wait until response accepted (r&v), then finish the miss
          lce_state_n = (lce_resp_ready_i) ? FINISH_MISS : LCE_CMD_STW_RESP;

        end
        FINISH_MISS: begin

          // send return packet back to TR after CCE handles the LCE miss request
          tr_pkt_v_o = 1'b1;
          tr_pkt_o[tr_ring_width_lp-1:dword_width_p] = '0;

          // TODO: return correct data for load
          tr_pkt_o[0 +: dword_width_p] = '0;
          if (load_op) begin
            // select data to return
            data_set = cmd.paddr[block_offset_bits_lp +: lg_lce_sets_lp];
            data_way = miss_lru_way_r;

            tr_pkt_o[0 +: dword_width_p] = double_op
              ? load_data
              : (word_op
                ? {{32{word_sigext}}, load_word}
                : (half_op
                  ? {{48{half_sigext}}, load_half}
                  : {{56{byte_sigext}}, load_byte}));
          end

          // wait until TR accepts packet (r&v), then go to READY
          if (tr_pkt_ready_i) begin
            lce_state_n = READY;

            // clear miss handling state
            miss_n = '0;
            miss_lru_way_n = '0;
            tag_received_n = '0;
            data_received_n = '0;

            // update lru_way
            lru_way_n = lru_way_r + 'd1;

          end else begin
            lce_state_n = FINISH_MISS;
          end

        end
        TR_CMD: begin
          // set up tag lookup
          tag_set = cmd.paddr[block_offset_bits_lp +: lg_lce_sets_lp];
          tag_set_li = tags[tag_set];
          ptag_li = cmd.paddr[paddr_width_p-1 -: ptag_width_lp];
          lru_way_li = lru_way_r;

          // tag_way depends on if there was a hit or not when it is a store
          tag_way = (tag_hit_lo) ? tag_hit_way_lo : '0;

          // capture tag lookup outputs
          tag_hit_n = tag_hit_lo;
          tag_dirty_n = tag_dirty_lo;
          tag_hit_way_n = tag_hit_way_lo;
          lru_dirty_n = lru_dirty_lo;

          // setup miss handling information
          miss_n = tag_hit_lo;
          miss_lru_way_n = lru_way_r;
          miss_st_upgrade_n = '0;
          tag_received_n = '0;
          data_received_n = '0;

          // process the trace replay command
          if (tag_hit_lo && load_op) begin
            lce_state_n = TR_CMD_LD_HIT;
          end else if (~tag_hit_lo && load_op) begin
            lce_state_n = TR_CMD_LD_MISS;
          end else if (~tag_hit_lo && store_op) begin
            lce_state_n = TR_CMD_ST_MISS;
          end else if (tag_hit_lo && store_op && ((tag_cur.coh_st == e_MESI_M) || (tag_cur.coh_st == e_MESI_E))) begin
            lce_state_n = TR_CMD_ST_HIT;
          end else if (tag_hit_lo && store_op && (tag_cur.coh_st == e_MESI_S)) begin
            miss_st_upgrade_n = 1'b1;
            lce_state_n = TR_CMD_ST_MISS;
          end else begin
            lce_state_n = RESET;
            $error("bad tag lookup");
          end

        end
        TR_CMD_LD_HIT: begin
          // load hit
          data_set = cmd.paddr[block_offset_bits_lp +: lg_lce_sets_lp];
          data_way = tag_hit_way_r;

          tr_pkt_v_o = 1'b1;
          tr_pkt_o[tr_ring_width_lp-1:dword_width_p] = '0;
          // select data to return
          tr_pkt_o[0 +: dword_width_p] = double_op
            ? load_data
            : (word_op
              ? {{32{word_sigext}}, load_word}
              : (half_op
                ? {{48{half_sigext}}, load_half}
                : {{56{byte_sigext}}, load_byte}));

          lce_state_n = (tr_pkt_ready_i) ? READY : TR_CMD_LD_HIT;

          // reset some state
          tag_hit_n = '0;
          tag_dirty_n = '0;
          tag_hit_way_n = '0;
          lru_dirty_n = '0;

          miss_n = '0;
          miss_lru_way_n = '0;
          miss_st_upgrade_n = '0;
          tag_received_n = '0;
          data_received_n = '0;

        end
        TR_CMD_LD_MISS: begin
          // load miss, send lce request
          lce_req_v_o = 1'b1;

          // TODO: in system with multiple CCE< dst_id needs to be computed from address
          lce_req_s.dst_id = '0;
          lce_req_s.src_id = lce_id_i;
          lce_req_s.data = '0;
          lce_req_s.msg_type = e_lce_req_type_rd;
          lce_req_s.non_exclusive = e_lce_req_excl;
          lce_req_s.addr = cmd.paddr;
          lce_req_s.lru_way_id = lru_way_r;
          lce_req_s.lru_dirty = (lru_dirty_r ? e_lce_req_lru_dirty : e_lce_req_lru_clean);
          lce_req_s.non_cacheable = e_lce_req_cacheable;
          lce_req_s.nc_size = e_lce_nc_req_1;

          // wait for LCE req outbound to be ready (r&v), then wait for responses
          lce_state_n = (lce_req_ready_i) ? READY : TR_CMD_LD_MISS;

        end
        TR_CMD_ST_HIT: begin
          // store hit on Exclusive forces upgrade to Modified
          tag_set = cmd.paddr[block_offset_bits_lp +: lg_lce_sets_lp];
          tag_way = tag_hit_way_r;
          if (tag_cur.coh_st == e_MESI_E) begin
            tag_w[tag_set][tag_way] = 1'b1;
            tag_n[tag_set][tag_way].coh_st = e_MESI_M;
            tag_n[tag_set][tag_way].tag = cmd.paddr[paddr_width_p-1 -: ptag_width_lp];
          end

          data_set = cmd.paddr[block_offset_bits_lp +: lg_lce_sets_lp];
          data_way = tag_hit_way_r;

          // TODO
          // do the store
          data_w[data_set][data_way] = 1'b1;
          data_mask_n = double_op
            ? {{(cce_block_width_p-64){1'b0}}, {64{1'b1}}} << (dword_offset*64)
            : word_op
              ? {{(cce_block_width_p-32){1'b0}}, {32{1'b1}}} << (dword_offset*64 + 32*byte_offset[2])
              : half_op
                ? {{(cce_block_width_p-16){1'b0}}, {16{1'b1}}} << (dword_offset*64 + 16*byte_offset[2:1])
                : {{(cce_block_width_p-8){1'b0}}, {8{1'b1}}} << (dword_offset*64 + 8*byte_offset[2:0]);

          data_n = double_op
            ? {{(cce_block_width_p-64){1'b0}}, cmd.data} << (dword_offset*64)
            : word_op
              ? {{(cce_block_width_p-32){1'b0}}, cmd.data[0+:32]} << (dword_offset*64 + 32*byte_offset[2])
              : half_op
                ? {{(cce_block_width_p-16){1'b0}}, cmd.data[0+:16]} << (dword_offset*64 + 16*byte_offset[2:1])
                : {{(cce_block_width_p-8){1'b0}}, cmd.data[0+:8]} << (dword_offset*64 + 8*byte_offset[2:0]);


          lce_state_n = TR_CMD_ST_HIT_RESP;
        end
        TR_CMD_ST_HIT_RESP: begin
          // reset some state
          tag_hit_n = '0;
          tag_dirty_n = '0;
          tag_hit_way_n = '0;
          lru_dirty_n = '0;

          miss_n = '0;
          miss_lru_way_n = '0;
          miss_st_upgrade_n = '0;
          tag_received_n = '0;
          data_received_n = '0;

          // output valid trace replay return packet
          tr_pkt_v_o = 1'b1;
          tr_pkt_o = '0;
          // wait until packet consumed, then go to ready
          lce_state_n = (tr_pkt_ready_i) ? READY : TR_CMD_ST_HIT_RESP;

        end
        TR_CMD_ST_MISS: begin
          // store miss - block present, not writable
          lce_req_v_o = 1'b1;

          lce_req_s.dst_id = '0;
          lce_req_s.src_id = lce_id_i;
          lce_req_s.data = '0;
          lce_req_s.msg_type = e_lce_req_type_wr;
          lce_req_s.non_exclusive = e_lce_req_excl;
          lce_req_s.addr = cmd.paddr;

          lce_req_s.lru_way_id = (miss_st_upgrade_r) ? tag_hit_way_r : miss_lru_way_r;
          lce_req_s.lru_dirty = (miss_st_upgrade_r) ? e_lce_req_lru_clean :
            ((lru_dirty_r) ? e_lce_req_lru_dirty : e_lce_req_lru_clean);
          
          lce_req_s.non_cacheable = e_lce_req_cacheable;
          lce_req_s.nc_size = e_lce_nc_req_1;

          lce_state_n = (lce_req_ready_i) ? READY : TR_CMD_ST_MISS;

        end
        default: begin
          lce_state_n = RESET;
        end
      endcase
    end
  end

  always_ff @(negedge clk_i) begin
      case (lce_state)
        TR_CMD: begin
          if (tag_hit_lo && load_op) begin
            $display("Load hit: M[%d]", cmd.paddr);
          end else if (~tag_hit_lo && load_op) begin
            $display("Load miss: M[%d]", cmd.paddr);
          end else if (~tag_hit_lo && store_op) begin
            $display("Store miss: M[%d] := %d", cmd.paddr, cmd.data);
          end else if (tag_hit_lo && store_op && ((tag_cur.coh_st == e_MESI_M) || (tag_cur.coh_st == e_MESI_E))) begin
            $display("Store hit: M[%d] := %d", cmd.paddr, cmd.data);
          end else if (tag_hit_lo && store_op && (tag_cur.coh_st == e_MESI_S)) begin
            $display("Store miss: M[%d] := %d", cmd.paddr, cmd.data);
          end
        end
      endcase

  end

endmodule


