/**
 *  Name:
 *    bp_me_wormhole_packet_encode_lce_cmd.v
 *
 *  Description:
 *    It takes bp_lce_cmd_s as a payload, parses, and forms it into a wormhole
 *    packet that goes into the adapter.
 *
 *    packet = {payload, length, cord}
 */


module bp_me_wormhole_packet_encode_lce_cmd
  import bp_common_pkg::*;
  import bp_common_aviary_pkg::*;
  #(parameter bp_cfg_e cfg_p = e_bp_inv_cfg
    `declare_bp_proc_params(cfg_p)
    `declare_bp_lce_cce_if_widths(num_cce_p, num_lce_p, paddr_width_p, lce_assoc_p, dword_width_p, cce_block_width_p)

    // Generalized Wormhole Router parameters
    , localparam dims_lp                                = 2
    , localparam coh_x_cord_width_lp                    = `BSG_SAFE_CLOG2(num_lce_p)
    , localparam coh_y_cord_width_lp                    = 1
    , localparam int coh_cord_markers_pos_lp[dims_lp:0] =
     '{ coh_x_cord_width_lp+coh_y_cord_width_lp, coh_x_cord_width_lp, 0 }
    , localparam coh_cord_width_lp = coh_cord_markers_pos_lp[dims_lp]

    , localparam lce_cmd_packet_width_lp = 
        `bsg_wormhole_concentrator_packet_width(coh_cord_width_lp, coh_noc_len_width_p, coh_noc_cid_width_p, lce_cmd_width_lp)
    )
   (input [lce_cmd_width_lp-1:0]           payload_i
    , output [lce_cmd_packet_width_lp-1:0] packet_o
    );

  `declare_bp_lce_cce_if(num_cce_p, num_lce_p, paddr_width_p, lce_assoc_p, dword_width_p, cce_block_width_p);
  `declare_bsg_wormhole_concentrator_packet_s(coh_cord_width_lp, coh_noc_len_width_p, coh_noc_cid_width_p, lce_cmd_width_lp, lce_cmd_packet_s);

  bp_lce_cmd_s payload_cast_i;
  lce_cmd_packet_s packet_cast_o;
  assign payload_cast_i = payload_i;
  assign packet_o = packet_cast_o;

  localparam lce_cmd_cmd_len_lp = 
    `BSG_CDIV(lce_cmd_packet_width_lp-$bits(payload_cast_i.msg.cmd.pad), coh_noc_flit_width_p) - 1;
  localparam lce_cmd_data_len_lp = 
    `BSG_CDIV(lce_cmd_packet_width_lp, coh_noc_flit_width_p) - 1;
  localparam lce_cmd_uc_data_len_lp =
    `BSG_CDIV(lce_cmd_packet_width_lp-(cce_block_width_p-dword_width_p), coh_noc_flit_width_p) - 1;

  always_comb begin
    packet_cast_o.payload = payload_cast_i;
    packet_cast_o.cid     = 1'b0;
    packet_cast_o.cord    = payload_cast_i.dst_id;

    case (payload_cast_i.msg_type)
      e_lce_cmd_sync
      ,e_lce_cmd_set_clear
      ,e_lce_cmd_transfer
      ,e_lce_cmd_writeback
      ,e_lce_cmd_set_tag
      ,e_lce_cmd_set_tag_wakeup
      ,e_lce_cmd_invalidate_tag
      ,e_lce_cmd_uc_st_done: packet_cast_o.len = lce_cmd_cmd_len_lp;
      e_lce_cmd_data       : packet_cast_o.len = lce_cmd_data_len_lp;
      e_lce_cmd_uc_data    : packet_cast_o.len = lce_cmd_uc_data_len_lp; 
      default: packet_cast_o = '0;
    endcase
  end

endmodule

