
package bp_fe_icache_pkg;

`include "bp_common_bedrock_if.vh"
`include "bsg_defines.v"
`include "bp_fe_icache.vh"

endpackage : bp_fe_icache_pkg
