
package bp_be_pkg;
  import bp_common_pkg::*;
  import bp_common_rv64_pkg::*;

  `include "bp_common_fe_be_if.vh"
  `include "bp_be_ctl_defines.vh"
  `include "bp_be_mem_defines.vh"
  `include "bp_be_internal_if_defines.vh"

endpackage : bp_be_pkg

