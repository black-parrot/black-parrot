`ifndef BP_TOP_DEFINES_SVH
`define BP_TOP_DEFINES_SVH

`endif

