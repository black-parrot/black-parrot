module wrapper
  import bp_common_pkg::*;
  import bp_common_aviary_pkg::*;
  import bp_common_cfg_link_pkg::*;
  import bp_fe_pkg::*;
  import bp_fe_icache_pkg::*;
  import bp_cce_pkg::*;
  import bp_me_pkg::*;
  #(parameter bp_params_e bp_params_p = BP_CFG_FLOWVAR
  `declare_bp_proc_params(bp_params_p)
  `declare_bp_fe_tag_widths(icache_assoc_p, lce_sets_p, lce_id_width_p, cce_id_width_p, dword_width_p, paddr_width_p)
  `declare_bp_cache_service_if_widths(paddr_width_p, ptag_width_p, lce_sets_p, icache_assoc_p, dword_width_p, cce_block_width_p, icache)
  `declare_bp_lce_cce_if_widths(cce_id_width_p, lce_id_width_p, paddr_width_p, lce_assoc_p, dword_width_p, cce_block_width_p)
  `declare_bp_me_if_widths(paddr_width_p, cce_block_width_p, lce_id_width_p, lce_assoc_p)

  , localparam cfg_bus_width_lp = `bp_cfg_bus_width(vaddr_width_p, core_id_width_p, cce_id_width_p, lce_id_width_p, cce_pc_width_p, cce_instr_width_p)
  , localparam lg_icache_assoc_lp = `BSG_SAFE_CLOG2(icache_assoc_p)
  , localparam way_id_width_lp=`BSG_SAFE_CLOG2(icache_assoc_p)
  , localparam block_size_in_words_lp=icache_assoc_p
  , localparam cache_block_width_multiplier_lp = 2**(3-`BSG_SAFE_CLOG2(icache_assoc_p))
  , localparam cache_block_width_lp = dword_width_p * cache_block_width_multiplier_lp
  , localparam data_mem_mask_width_lp=(cache_block_width_lp>>3)
  , localparam byte_offset_width_lp=`BSG_SAFE_CLOG2(cache_block_width_lp>>3)
  , localparam word_offset_width_lp=`BSG_SAFE_CLOG2(block_size_in_words_lp)
  , localparam index_width_lp=`BSG_SAFE_CLOG2(lce_sets_p)
  , localparam block_offset_width_lp=(word_offset_width_lp+byte_offset_width_lp)
  , localparam ptag_width_lp=(paddr_width_p-bp_page_offset_width_gp)
  , localparam stat_width_lp = `bp_be_dcache_stat_info_width(icache_assoc_p) 
 
  )
  ( input                             clk_i
  , input                             reset_i

  , input [cfg_bus_width_lp-1:0]      cfg_bus_i

  , input [vaddr_width_p-1:0]         vaddr_i
  , input                             vaddr_v_i
  , input                             fencei_v_i
  , output                            vaddr_ready_o

  , input [ptag_width_p-1:0]          ptag_i
  , input                             ptag_v_i
  , input                             uncached_i
  , input                             poison_i

  , output [instr_width_p-1:0]        data_o
  , output                            data_v_o
  , output                            miss_o

  , input [cce_mem_msg_width_lp-1:0]  mem_resp_i
  , input                             mem_resp_v_i
  , output                            mem_resp_ready_o

  , output [cce_mem_msg_width_lp-1:0] mem_cmd_o
  , output                            mem_cmd_v_o
  , input                             mem_cmd_yumi_i
  );

  // I$-LCE Interface signals
  // Miss, Management Interfaces
  logic cache_req_ready_li;
  logic [cache_req_width_lp-1:0] cache_req_lo;
  logic cache_req_v_lo;
  logic [cache_req_metadata_width_lp-1:0] cache_req_metadata_lo;
  logic cache_req_metadata_v_lo;

  logic cache_req_complete_li;

  // Fill Interfaces
  logic data_mem_pkt_v_li, tag_mem_pkt_v_li, stat_mem_pkt_v_li;
  logic data_mem_pkt_ready_lo, tag_mem_pkt_ready_lo, stat_mem_pkt_ready_lo;
  logic [icache_data_mem_pkt_width_lp-1:0] data_mem_pkt_li;
  logic [icache_tag_mem_pkt_width_lp-1:0] tag_mem_pkt_li;
  logic [icache_stat_mem_pkt_width_lp-1:0] stat_mem_pkt_li;
  logic [cce_block_width_p-1:0] data_mem_lo;
  logic [ptag_width_lp-1:0] tag_mem_lo;
  logic [stat_width_lp-1:0] stat_mem_lo;
  
  // LCE-CCE Interface
  logic lce_req_v_lo, lce_resp_v_lo, lce_cmd_v_li;
  logic lce_req_ready_li, lce_resp_ready_li, lce_cmd_yumi_lo;
  logic [lce_cce_req_width_lp-1:0] lce_req_lo;
  logic [lce_cce_resp_width_lp-1:0] lce_resp_lo;
  logic [lce_cmd_width_lp-1:0] lce_cmd_li;

  // TODO: Add a rolly fifo here

  // I-Cache
  bp_fe_icache
    #(.bp_params_p(bp_params_p))
    icache
    (.clk_i(clk_i)
    ,.reset_i(reset_i)
    
    ,.cfg_bus_i(cfg_bus_i)
    
    ,.vaddr_i(vaddr_i)
    ,.vaddr_v_i(vaddr_v_i)
    ,.fencei_v_i(fencei_v_i)
    ,.vaddr_ready_o(vaddr_ready_o)    

    ,.ptag_i(ptag_i)
    ,.ptag_v_i(ptag_v_i)
    ,.uncached_i(uncached_i)
    ,.poison_i(poison_i)

    ,.data_o(data_o)
    ,.data_v_o(data_v_o)
    ,.miss_o(miss_o)
     
    ,.cache_req_ready_i(cache_req_ready_li)
    ,.cache_req_o(cache_req_lo)
    ,.cache_req_v_o(cache_req_v_lo)
    ,.cache_req_metadata_o(cache_req_metadata_lo)
    ,.cache_req_metadata_v_o(cache_req_metadata_v_lo)

    ,.cache_req_complete_i(cache_req_complete_li)

    ,.data_mem_pkt_v_i(data_mem_pkt_v_li)
    ,.data_mem_pkt_i(data_mem_pkt_li)
    ,.data_mem_o(data_mem_lo)
    ,.data_mem_pkt_ready_o(data_mem_pkt_ready_lo)

    ,.tag_mem_pkt_v_i(tag_mem_pkt_v_li)
    ,.tag_mem_pkt_i(tag_mem_pkt_li)
    ,.tag_mem_o(tag_mem_lo)
    ,.tag_mem_pkt_ready_o(tag_mem_pkt_ready_lo)

    ,.stat_mem_pkt_v_i(stat_mem_pkt_v_li)
    ,.stat_mem_pkt_i(stat_mem_pkt_li)
    ,.stat_mem_o(stat_mem_lo)
    ,.stat_mem_pkt_ready_o(stat_mem_pkt_ready_lo)
    );

  // I-Cache LCE
  bp_fe_lce
    #(.bp_params_p(bp_params_p))
    icache_lce
    (.clk_i(clk_i)
    ,.reset_i(reset_i)
    
    ,.cfg_bus_i(cfg_bus_i)

    ,.cache_req_v_i(cache_req_v_lo)
    ,.cache_req_i(cache_req_lo)
    ,.cache_req_ready_o(cache_req_ready_li)
    ,.cache_req_metadata_i(cache_req_metadata_lo)
    ,.cache_req_metadata_v_i(cache_req_metadata_v_lo)

    ,.cache_req_complete_o(cache_req_complete_li)

    ,.data_mem_i(data_mem_lo)
    ,.data_mem_pkt_o(data_mem_pkt_li)
    ,.data_mem_pkt_v_o(data_mem_pkt_v_li)
    ,.data_mem_pkt_ready_i(data_mem_pkt_ready_lo)
    
    ,.tag_mem_i(tag_mem_lo)
    ,.tag_mem_pkt_o(tag_mem_pkt_li)
    ,.tag_mem_pkt_v_o(tag_mem_pkt_v_li)
    ,.tag_mem_pkt_ready_i(tag_mem_pkt_ready_lo)

    ,.stat_mem_i(stat_mem_lo)
    ,.stat_mem_pkt_o(stat_mem_pkt_li)
    ,.stat_mem_pkt_v_o(stat_mem_pkt_v_li)
    ,.stat_mem_pkt_ready_i(stat_mem_pkt_ready_lo)

    ,.lce_req_o(lce_req_lo)
    ,.lce_req_v_o(lce_req_v_lo)
    ,.lce_req_ready_i(lce_req_ready_li)

    ,.lce_resp_o(lce_resp_lo)
    ,.lce_resp_v_o(lce_resp_v_lo)
    ,.lce_resp_ready_i(lce_resp_ready_li)

    ,.lce_cmd_i(lce_cmd_li)
    ,.lce_cmd_v_i(lce_cmd_v_li)
    ,.lce_cmd_yumi_o(lce_cmd_yumi_lo)

    ,.lce_cmd_o()
    ,.lce_cmd_v_o()
    ,.lce_cmd_ready_i()
    );  
 
  bp_cce_fsm_top
  	#(.bp_params_p(bp_params_p))
  	cce_top
  	(.clk_i(clk_i)
  	,.reset_i(reset_i)

  	,.cfg_bus_i(cfg_bus_i)
  	,.cfg_cce_ucode_data_o()

  	,.lce_req_i(lce_req_lo)
  	,.lce_req_v_i(lce_req_v_lo)
  	,.lce_req_ready_o(lce_req_ready_li)

  	,.lce_resp_i(lce_resp_lo)
  	,.lce_resp_v_i(lce_resp_v_lo)
  	,.lce_resp_ready_o(lce_resp_ready_li)

  	,.lce_cmd_o(lce_cmd_li)
  	,.lce_cmd_v_o(lce_cmd_v_li)
  	,.lce_cmd_ready_i(lce_cmd_yumi_lo)

  	,.mem_resp_i(mem_resp_i)
  	,.mem_resp_v_i(mem_resp_v_i)
  	,.mem_resp_ready_o(mem_resp_ready_o)

  	,.mem_cmd_o(mem_cmd_o)
  	,.mem_cmd_v_o(mem_cmd_v_o)
  	,.mem_cmd_yumi_i(mem_cmd_yumi_i)
  	); 

endmodule  
